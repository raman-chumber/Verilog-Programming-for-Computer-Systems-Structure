//4x1 Multiplexer by Ramandeep Chumber
 module MuxMod(s1, s0, d0, d1, d2, d3, o);
input s1, s0, d0, d1, d2, d3;
   output o;

   wire s1_inv, s0_inv, and0, and1, and2, and3, and4, and5, and6, and7, or0, or1;

   not(s1_inv, s1);
   not(s0_inv, s0);

   and(and0, d0, s1_inv);
   and(and1, and0, s0_inv);

   and(and2, d1, s1_inv);
   and(and3, and2, s0);

   and(and4, d2, s1);
   and(and5, and4, s0_inv);

   and(and6, d3, s1);
   and(and7, and6, s0);

   or(or0, and1, and3);      // "or" is a built-in gate
   or(or1, and5, and7);      // "or" is a built-in gate

   or(o, or0, or1);      // "or" is a built-in gate
endmodule

module TestMod;
   reg s1, s0, d0, d1, d2, d3;
   wire o;

   MuxMod my_mux(s1, s0, d0, d1, d2, d3, o);
    initial begin
      $display("Time s1 s0 d0 d1 d2 d3  o");
      $display("-------------------------");
      $monitor("%3d   %b  %b  %b  %b  %b  %b  %b",
         $time, s1, s0, d0, d1, d2, d3, o);
   end

   initial #63 $finish;

   initial begin
            s1=0; s0=0; d0=0; d1=0; d2=0; d3=0;
      #1 s1=0; s0=0; d0=0; d1=0; d2=0; d3=1;
      #1 s1=0; s0=0; d0=0; d1=0; d2=1; d3=0;
      #1 s1=0; s0=0; d0=0; d1=0; d2=1; d3=1;
      #1 s1=0; s0=0; d0=0; d1=1; d2=0; d3=0;
      #1 s1=0; s0=0; d0=0; d1=1; d2=0; d3=1;
      #1 s1=0; s0=0; d0=0; d1=1; d2=1; d3=0;
      #1 s1=0; s0=0; d0=0; d1=1; d2=1; d3=1;
      #1 s1=0; s0=0; d0=1; d1=0; d2=0; d3=0;
      #1 s1=0; s0=0; d0=1; d1=0; d2=0; d3=1;
      #1 s1=0; s0=0; d0=1; d1=0; d2=1; d3=0;
      #1 s1=0; s0=0; d0=1; d1=0; d2=1; d3=1;
      #1 s1=0; s0=0; d0=1; d1=1; d2=0; d3=0;
      #1 s1=0; s0=0; d0=1; d1=1; d2=0; d3=1;
      #1 s1=0; s0=0; d0=1; d1=1; d2=1; d3=0;
      #1 s1=0; s0=0; d0=1; d1=1; d2=1; d3=1;
      #1 s1=0; s0=1; d0=0; d1=0; d2=0; d3=0;
      #1 s1=0; s0=1; d0=0; d1=0; d2=0; d3=1;
      #1 s1=0; s0=1; d0=0; d1=0; d2=1; d3=0;
      #1 s1=0; s0=1; d0=0; d1=0; d2=1; d3=1;
      #1 s1=0; s0=1; d0=0; d1=1; d2=0; d3=0;
      #1 s1=0; s0=1; d0=0; d1=1; d2=0; d3=1;
      #1 s1=0; s0=1; d0=0; d1=1; d2=1; d3=0;
      #1 s1=0; s0=1; d0=0; d1=1; d2=1; d3=1;
      #1 s1=0; s0=1; d0=1; d1=0; d2=0; d3=0;
      #1 s1=0; s0=1; d0=1; d1=0; d2=0; d3=1;
      #1 s1=0; s0=1; d0=1; d1=0; d2=1; d3=0;
      #1 s1=0; s0=1; d0=1; d1=0; d2=1; d3=1;
      #1 s1=0; s0=1; d0=1; d1=1; d2=0; d3=0;
      #1 s1=0; s0=1; d0=1; d1=1; d2=0; d3=1;
      #1 s1=0; s0=1; d0=1; d1=1; d2=1; d3=0;
      #1 s1=0; s0=1; d0=1; d1=1; d2=1; d3=1;
      #1 s1=1; s0=0; d0=0; d1=0; d2=0; d3=0;
      #1 s1=1; s0=0; d0=0; d1=0; d2=0; d3=1;
      #1 s1=1; s0=0; d0=0; d1=0; d2=1; d3=0;
      #1 s1=1; s0=0; d0=0; d1=0; d2=1; d3=1;
      #1 s1=1; s0=0; d0=0; d1=1; d2=0; d3=0;
      #1 s1=1; s0=0; d0=0; d1=1; d2=0; d3=1;
      #1 s1=1; s0=0; d0=0; d1=1; d2=1; d3=0;
      #1 s1=1; s0=0; d0=0; d1=1; d2=1; d3=1;
      #1 s1=1; s0=0; d0=1; d1=0; d2=0; d3=0;
      #1 s1=1; s0=0; d0=1; d1=0; d2=0; d3=1;
      #1 s1=1; s0=0; d0=1; d1=0; d2=1; d3=0;
      #1 s1=1; s0=0; d0=1; d1=0; d2=1; d3=1;
      #1 s1=1; s0=0; d0=1; d1=1; d2=0; d3=0;
      #1 s1=1; s0=0; d0=1; d1=1; d2=0; d3=1;
      #1 s1=1; s0=0; d0=1; d1=1; d2=1; d3=0;
      #1 s1=1; s0=0; d0=1; d1=1; d2=1; d3=1;
      #1 s1=1; s0=1; d0=0; d1=0; d2=0; d3=0;
      #1 s1=1; s0=1; d0=0; d1=0; d2=0; d3=1;
      #1 s1=1; s0=1; d0=0; d1=0; d2=1; d3=0;
      #1 s1=1; s0=1; d0=0; d1=0; d2=1; d3=1;
      #1 s1=1; s0=1; d0=0; d1=1; d2=0; d3=0;
      #1 s1=1; s0=1; d0=0; d1=1; d2=0; d3=1;
      #1 s1=1; s0=1; d0=0; d1=1; d2=1; d3=0;
      #1 s1=1; s0=1; d0=0; d1=1; d2=1; d3=1;
      #1 s1=1; s0=1; d0=1; d1=0; d2=0; d3=0;
      #1 s1=1; s0=1; d0=1; d1=0; d2=0; d3=1;
      #1 s1=1; s0=1; d0=1; d1=0; d2=1; d3=0;
      #1 s1=1; s0=1; d0=1; d1=0; d2=1; d3=1;
      #1 s1=1; s0=1; d0=1; d1=1; d2=0; d3=0;
      #1 s1=1; s0=1; d0=1; d1=1; d2=0; d3=1;
      #1 s1=1; s0=1; d0=1; d1=1; d2=1; d3=0;
      #1 s1=1; s0=1; d0=1; d1=1; d2=1; d3=1;
   end
endmodule